module sorting_box#(
    parameter DATA_WD = 8,
    parameter SIGNED=0
)(
    input   logic   [DATA_WD-1:0]   i_a[4],
    output  logic   [DATA_WD-1:0]   o_sorted_a[4]
);


endmodule
